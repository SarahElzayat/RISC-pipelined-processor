module processor(
    input clk,
    input rst
);

endmodule 
