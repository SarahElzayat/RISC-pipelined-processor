module name(
    input clk,
    input rst
);
    
endmodule : name
